//
// This module synchronizes, debounces, and one-pulses a button input.
//
module button_process_unit(
  input clk,
  input reset,
  input ButtonIn,
  output ButtonOut
  );
  
endmodule
   